`ifndef TYPES
`define TYPES


localparam int gRegs        = 16;
localparam int gDataWidth   = 16;

typedef bit[gDataWidth-1 : 0] data_v;


`endif
