`ifndef TYPES
`define TYPES


localparam int gRegs = 16;

typedef bit[gRegs-1 : 0] data_v;


`endif
