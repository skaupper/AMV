`ifndef _CHECKER_
`define _CHECKER_

`include "types.sv"

class Checker;


endclass


`endif /* _CHECKER_ */
