`ifndef _DRIVER_
`define _DRIVER_

`include "types.sv"

class Driver;


endclass


`endif /* _DRIVER_ */
