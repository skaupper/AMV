entity WishboneBFM_tb is
end entity;

architecture tb of WishboneBFM_tb is

begin



end architecture tb;
