`ifndef _DRIVER_
`define _DRIVER_

//`include

class Driver;


endclass


`endif /* _DRIVER_ */
