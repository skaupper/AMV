`ifndef _AGENT_
`define _AGENT_

`include "types.sv"

class Agent;


endclass


`endif /* _AGENT_ */
