package WishboneBFM_pack is
end package;

package body WishboneBFM_pack is

end package body;
